library IEEE;
use IEEE.std_logic_1164.all;

entity pipeline is
	port( CLK	: in std_logic);
end pipeline;

architecture BV of pipeline is










end BV;